-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity coco3_Char_ROM is
  port (
    CLK         : in    std_logic;
    ADDR_R      : in    std_logic_vector(11 downto 0);
    ADDR_W      : in    std_logic_vector(11 downto 0);
	WE			: in    std_logic;
    DATA_R      : out   std_logic_vector(7 downto 0);
    DATA_W      : in    std_logic_vector(7 downto 0)
    );
end;

architecture RTL of coco3_Char_ROM is


  type RAM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  signal RAM : RAM_ARRAY := (
    x"00",x"00",x"00",x"1C",x"22",x"20",x"20",x"20", -- 0x0000
    x"22",x"1C",x"08",x"00",x"00",x"00",x"00",x"00", -- 0x0008
    x"00",x"00",x"00",x"22",x"00",x"22",x"22",x"22", -- 0x0010
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0018
    x"00",x"00",x"00",x"04",x"08",x"1C",x"22",x"3E", -- 0x0020
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0028
    x"00",x"00",x"00",x"08",x"14",x"1C",x"02",x"1E", -- 0x0030
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0038
    x"00",x"00",x"00",x"14",x"00",x"1C",x"02",x"1E", -- 0x0040
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0048
    x"00",x"00",x"00",x"10",x"08",x"1C",x"02",x"1E", -- 0x0050
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"08",x"00",x"1C",x"02",x"1E", -- 0x0060
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0068
    x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"20", -- 0x0070
    x"22",x"1C",x"08",x"00",x"00",x"00",x"00",x"00", -- 0x0078
    x"00",x"00",x"00",x"08",x"14",x"1C",x"22",x"3E", -- 0x0080
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0088
    x"00",x"00",x"00",x"14",x"00",x"1C",x"22",x"3E", -- 0x0090
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0098
    x"00",x"00",x"00",x"10",x"08",x"1C",x"22",x"3E", -- 0x00A0
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A8
    x"00",x"00",x"00",x"14",x"00",x"18",x"08",x"08", -- 0x00B0
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B8
    x"00",x"00",x"00",x"08",x"14",x"00",x"18",x"08", -- 0x00C0
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C8
    x"00",x"00",x"00",x"00",x"0C",x"12",x"1C",x"12", -- 0x00D0
    x"12",x"1C",x"20",x"00",x"00",x"00",x"00",x"00", -- 0x00D8
    x"00",x"00",x"00",x"22",x"08",x"14",x"22",x"3E", -- 0x00E0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E8
    x"00",x"00",x"00",x"08",x"08",x"14",x"22",x"3E", -- 0x00F0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F8
    x"00",x"00",x"00",x"04",x"08",x"1C",x"22",x"22", -- 0x0100
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0108
    x"00",x"00",x"00",x"00",x"00",x"34",x"0A",x"1E", -- 0x0110
    x"28",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0118
    x"00",x"00",x"00",x"1E",x"28",x"28",x"3C",x"28", -- 0x0120
    x"28",x"2C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0128
    x"00",x"00",x"00",x"08",x"14",x"1C",x"22",x"22", -- 0x0130
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0138
    x"00",x"00",x"00",x"14",x"00",x"1C",x"22",x"22", -- 0x0140
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0148
    x"00",x"00",x"00",x"00",x"00",x"1C",x"26",x"2E", -- 0x0150
    x"32",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0158
    x"00",x"00",x"00",x"08",x"14",x"00",x"22",x"22", -- 0x0160
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0168
    x"00",x"00",x"00",x"10",x"08",x"22",x"22",x"22", -- 0x0170
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"00",x"1C",x"26",x"2A",x"2A",x"2A", -- 0x0180
    x"32",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0188
    x"00",x"00",x"00",x"22",x"1C",x"22",x"22",x"22", -- 0x0190
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"14",x"22",x"22",x"22",x"22", -- 0x01A0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
    x"00",x"00",x"00",x"1C",x"20",x"1C",x"22",x"1C", -- 0x01B0
    x"02",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
    x"00",x"00",x"00",x"04",x"0A",x"08",x"1C",x"08", -- 0x01C0
    x"0A",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
    x"00",x"00",x"00",x"08",x"08",x"3E",x"08",x"08", -- 0x01D0
    x"00",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D8
    x"00",x"00",x"00",x"04",x"0A",x"04",x"00",x"00", -- 0x01E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
    x"00",x"00",x"00",x"04",x"0A",x"08",x"1C",x"08", -- 0x01F0
    x"08",x"28",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0208
    x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"08", -- 0x0210
    x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0218
    x"00",x"00",x"00",x"14",x"14",x"14",x"00",x"00", -- 0x0220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0228
    x"00",x"00",x"00",x"14",x"14",x"3E",x"14",x"3E", -- 0x0230
    x"14",x"14",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0238
    x"00",x"00",x"00",x"08",x"1E",x"28",x"1C",x"0A", -- 0x0240
    x"3C",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0248
    x"00",x"00",x"00",x"32",x"32",x"04",x"08",x"10", -- 0x0250
    x"26",x"26",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0258
    x"00",x"00",x"00",x"10",x"28",x"28",x"10",x"2A", -- 0x0260
    x"24",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
    x"00",x"00",x"00",x"08",x"08",x"10",x"00",x"00", -- 0x0270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0278
    x"00",x"00",x"00",x"08",x"10",x"20",x"20",x"20", -- 0x0280
    x"10",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
    x"00",x"00",x"00",x"08",x"04",x"02",x"02",x"02", -- 0x0290
    x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0298
    x"00",x"00",x"00",x"00",x"08",x"2A",x"1C",x"1C", -- 0x02A0
    x"2A",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
    x"00",x"00",x"00",x"00",x"08",x"08",x"3E",x"08", -- 0x02B0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C0
    x"08",x"08",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x02C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"00", -- 0x02D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E0
    x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E8
    x"00",x"00",x"00",x"00",x"02",x"04",x"08",x"10", -- 0x02F0
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"00",x"00",x"00",x"1C",x"22",x"26",x"2A",x"32", -- 0x0300
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0308
    x"00",x"00",x"00",x"08",x"18",x"08",x"08",x"08", -- 0x0310
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0318
    x"00",x"00",x"00",x"1C",x"22",x"02",x"1C",x"20", -- 0x0320
    x"20",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0328
    x"00",x"00",x"00",x"1C",x"22",x"02",x"04",x"02", -- 0x0330
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0338
    x"00",x"00",x"00",x"04",x"0C",x"14",x"24",x"3E", -- 0x0340
    x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0348
    x"00",x"00",x"00",x"3E",x"20",x"3C",x"02",x"02", -- 0x0350
    x"02",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0358
    x"00",x"00",x"00",x"1C",x"20",x"20",x"3C",x"22", -- 0x0360
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0368
    x"00",x"00",x"00",x"3E",x"02",x"04",x"08",x"10", -- 0x0370
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0378
    x"00",x"00",x"00",x"1C",x"22",x"22",x"1C",x"22", -- 0x0380
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0388
    x"00",x"00",x"00",x"1C",x"22",x"22",x"1E",x"02", -- 0x0390
    x"02",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00", -- 0x03A0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
    x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00", -- 0x03B0
    x"08",x"08",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"04",x"08",x"10",x"20",x"10", -- 0x03C0
    x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"00",x"00",x"00",x"3E",x"00",x"3E", -- 0x03D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"00",x"00",x"00",x"10",x"08",x"04",x"02",x"04", -- 0x03E0
    x"08",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
    x"00",x"00",x"00",x"1C",x"22",x"02",x"04",x"08", -- 0x03F0
    x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
    x"00",x"00",x"00",x"1C",x"22",x"02",x"1A",x"2A", -- 0x0400
    x"2A",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0408
    x"00",x"00",x"00",x"08",x"14",x"22",x"22",x"3E", -- 0x0410
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0418
    x"00",x"00",x"00",x"3C",x"12",x"12",x"1C",x"12", -- 0x0420
    x"12",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0428
    x"00",x"00",x"00",x"1C",x"22",x"20",x"20",x"20", -- 0x0430
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
    x"00",x"00",x"00",x"3C",x"12",x"12",x"12",x"12", -- 0x0440
    x"12",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0448
    x"00",x"00",x"00",x"3E",x"20",x"20",x"3C",x"20", -- 0x0450
    x"20",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0458
    x"00",x"00",x"00",x"3E",x"20",x"20",x"3C",x"20", -- 0x0460
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0468
    x"00",x"00",x"00",x"1E",x"20",x"20",x"26",x"22", -- 0x0470
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0478
    x"00",x"00",x"00",x"22",x"22",x"22",x"3E",x"22", -- 0x0480
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0488
    x"00",x"00",x"00",x"1C",x"08",x"08",x"08",x"08", -- 0x0490
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0498
    x"00",x"00",x"00",x"02",x"02",x"02",x"02",x"22", -- 0x04A0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04A8
    x"00",x"00",x"00",x"22",x"24",x"28",x"30",x"28", -- 0x04B0
    x"24",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B8
    x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20", -- 0x04C0
    x"20",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04C8
    x"00",x"00",x"00",x"22",x"36",x"2A",x"2A",x"22", -- 0x04D0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04D8
    x"00",x"00",x"00",x"22",x"32",x"2A",x"26",x"22", -- 0x04E0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E8
    x"00",x"00",x"00",x"1C",x"22",x"22",x"22",x"22", -- 0x04F0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F8
    x"00",x"00",x"00",x"3C",x"22",x"22",x"3C",x"20", -- 0x0500
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0508
    x"00",x"00",x"00",x"1C",x"22",x"22",x"22",x"2A", -- 0x0510
    x"24",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0518
    x"00",x"00",x"00",x"3C",x"22",x"22",x"3C",x"28", -- 0x0520
    x"24",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0528
    x"00",x"00",x"00",x"1C",x"22",x"10",x"08",x"04", -- 0x0530
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0538
    x"00",x"00",x"00",x"3E",x"08",x"08",x"08",x"08", -- 0x0540
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0548
    x"00",x"00",x"00",x"22",x"22",x"22",x"22",x"22", -- 0x0550
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0558
    x"00",x"00",x"00",x"22",x"22",x"22",x"14",x"14", -- 0x0560
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0568
    x"00",x"00",x"00",x"22",x"22",x"22",x"2A",x"2A", -- 0x0570
    x"36",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0578
    x"00",x"00",x"00",x"22",x"22",x"14",x"08",x"14", -- 0x0580
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0588
    x"00",x"00",x"00",x"22",x"22",x"14",x"08",x"08", -- 0x0590
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0598
    x"00",x"00",x"00",x"3E",x"02",x"04",x"08",x"10", -- 0x05A0
    x"20",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A8
    x"00",x"00",x"00",x"38",x"20",x"20",x"20",x"20", -- 0x05B0
    x"20",x"38",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B8
    x"00",x"00",x"00",x"20",x"20",x"10",x"08",x"04", -- 0x05C0
    x"02",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C8
    x"00",x"00",x"00",x"0E",x"02",x"02",x"02",x"02", -- 0x05D0
    x"02",x"0E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D8
    x"00",x"00",x"00",x"08",x"1C",x"2A",x"08",x"08", -- 0x05E0
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E8
    x"00",x"00",x"00",x"00",x"08",x"10",x"3E",x"10", -- 0x05F0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F8
    x"00",x"00",x"00",x"08",x"14",x"22",x"00",x"00", -- 0x0600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0608
    x"00",x"00",x"00",x"00",x"00",x"1C",x"02",x"1E", -- 0x0610
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0618
    x"00",x"00",x"00",x"20",x"20",x"2C",x"32",x"22", -- 0x0620
    x"32",x"2C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0628
    x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"20", -- 0x0630
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0638
    x"00",x"00",x"00",x"02",x"02",x"1A",x"26",x"22", -- 0x0640
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0648
    x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"3E", -- 0x0650
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0658
    x"00",x"00",x"00",x"04",x"0A",x"08",x"1C",x"08", -- 0x0660
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0668
    x"00",x"00",x"00",x"00",x"00",x"1A",x"26",x"26", -- 0x0670
    x"1A",x"02",x"1C",x"00",x"00",x"00",x"00",x"00", -- 0x0678
    x"00",x"00",x"00",x"20",x"20",x"2C",x"32",x"22", -- 0x0680
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0688
    x"00",x"00",x"00",x"00",x"08",x"00",x"18",x"08", -- 0x0690
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0698
    x"00",x"00",x"00",x"00",x"02",x"00",x"02",x"02", -- 0x06A0
    x"02",x"22",x"1C",x"00",x"00",x"00",x"00",x"00", -- 0x06A8
    x"00",x"00",x"00",x"20",x"20",x"24",x"28",x"30", -- 0x06B0
    x"28",x"24",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06B8
    x"00",x"00",x"00",x"18",x"08",x"08",x"08",x"08", -- 0x06C0
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C8
    x"00",x"00",x"00",x"00",x"00",x"14",x"2A",x"2A", -- 0x06D0
    x"2A",x"2A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D8
    x"00",x"00",x"00",x"00",x"00",x"2C",x"32",x"22", -- 0x06E0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06E8
    x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"22", -- 0x06F0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06F8
    x"00",x"00",x"00",x"00",x"00",x"2C",x"32",x"32", -- 0x0700
    x"2C",x"20",x"20",x"00",x"00",x"00",x"00",x"00", -- 0x0708
    x"00",x"00",x"00",x"00",x"00",x"1A",x"26",x"26", -- 0x0710
    x"1A",x"02",x"02",x"00",x"00",x"00",x"00",x"00", -- 0x0718
    x"00",x"00",x"00",x"00",x"00",x"2C",x"32",x"20", -- 0x0720
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0728
    x"00",x"00",x"00",x"00",x"00",x"1E",x"20",x"1C", -- 0x0730
    x"02",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0738
    x"00",x"00",x"00",x"10",x"10",x"38",x"10",x"10", -- 0x0740
    x"12",x"0C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0748
    x"00",x"00",x"00",x"00",x"00",x"22",x"22",x"22", -- 0x0750
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0758
    x"00",x"00",x"00",x"00",x"00",x"22",x"22",x"22", -- 0x0760
    x"14",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0768
    x"00",x"00",x"00",x"00",x"00",x"22",x"2A",x"2A", -- 0x0770
    x"14",x"14",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
    x"00",x"00",x"00",x"00",x"00",x"22",x"14",x"08", -- 0x0780
    x"14",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0788
    x"00",x"00",x"00",x"00",x"00",x"22",x"22",x"22", -- 0x0790
    x"1E",x"02",x"1C",x"00",x"00",x"00",x"00",x"00", -- 0x0798
    x"00",x"00",x"00",x"00",x"00",x"3E",x"04",x"08", -- 0x07A0
    x"10",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A8
    x"00",x"00",x"00",x"08",x"10",x"10",x"20",x"10", -- 0x07B0
    x"10",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B8
    x"00",x"00",x"00",x"08",x"08",x"08",x"00",x"08", -- 0x07C0
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
    x"00",x"00",x"00",x"08",x"04",x"04",x"02",x"04", -- 0x07D0
    x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D8
    x"00",x"00",x"00",x"10",x"2A",x"04",x"00",x"00", -- 0x07E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F0
    x"00",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F8
	
    x"00",x"00",x"00",x"1C",x"22",x"20",x"20",x"20", -- 0x0000
    x"22",x"1C",x"08",x"00",x"00",x"00",x"00",x"00", -- 0x0008
    x"00",x"00",x"00",x"22",x"00",x"22",x"22",x"22", -- 0x0010
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0018
    x"00",x"00",x"00",x"04",x"08",x"1C",x"22",x"3E", -- 0x0020
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0028
    x"00",x"00",x"00",x"08",x"14",x"1C",x"02",x"1E", -- 0x0030
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0038
    x"00",x"00",x"00",x"14",x"00",x"1C",x"02",x"1E", -- 0x0040
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0048
    x"00",x"00",x"00",x"10",x"08",x"1C",x"02",x"1E", -- 0x0050
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"08",x"00",x"1C",x"02",x"1E", -- 0x0060
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0068
    x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"20", -- 0x0070
    x"22",x"1C",x"08",x"00",x"00",x"00",x"00",x"00", -- 0x0078
    x"00",x"00",x"00",x"08",x"14",x"1C",x"22",x"3E", -- 0x0080
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0088
    x"00",x"00",x"00",x"14",x"00",x"1C",x"22",x"3E", -- 0x0090
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0098
    x"00",x"00",x"00",x"10",x"08",x"1C",x"22",x"3E", -- 0x00A0
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A8
    x"00",x"00",x"00",x"14",x"00",x"18",x"08",x"08", -- 0x00B0
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B8
    x"00",x"00",x"00",x"08",x"14",x"00",x"18",x"08", -- 0x00C0
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C8
    x"00",x"00",x"00",x"00",x"0C",x"12",x"1C",x"12", -- 0x00D0
    x"12",x"1C",x"20",x"00",x"00",x"00",x"00",x"00", -- 0x00D8
    x"00",x"00",x"00",x"22",x"08",x"14",x"22",x"3E", -- 0x00E0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E8
    x"00",x"00",x"00",x"08",x"08",x"14",x"22",x"3E", -- 0x00F0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F8
    x"00",x"00",x"00",x"04",x"08",x"1C",x"22",x"22", -- 0x0100
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0108
    x"00",x"00",x"00",x"00",x"00",x"34",x"0A",x"1E", -- 0x0110
    x"28",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0118
    x"00",x"00",x"00",x"1E",x"28",x"28",x"3C",x"28", -- 0x0120
    x"28",x"2C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0128
    x"00",x"00",x"00",x"08",x"14",x"1C",x"22",x"22", -- 0x0130
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0138
    x"00",x"00",x"00",x"14",x"00",x"1C",x"22",x"22", -- 0x0140
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0148
    x"00",x"00",x"00",x"00",x"00",x"1C",x"26",x"2E", -- 0x0150
    x"32",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0158
    x"00",x"00",x"00",x"08",x"14",x"00",x"22",x"22", -- 0x0160
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0168
    x"00",x"00",x"00",x"10",x"08",x"22",x"22",x"22", -- 0x0170
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"00",x"1C",x"26",x"2A",x"2A",x"2A", -- 0x0180
    x"32",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0188
    x"00",x"00",x"00",x"22",x"1C",x"22",x"22",x"22", -- 0x0190
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"14",x"22",x"22",x"22",x"22", -- 0x01A0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
    x"00",x"00",x"00",x"1C",x"20",x"1C",x"22",x"1C", -- 0x01B0
    x"02",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
    x"00",x"00",x"00",x"04",x"0A",x"08",x"1C",x"08", -- 0x01C0
    x"0A",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
    x"00",x"00",x"00",x"08",x"08",x"3E",x"08",x"08", -- 0x01D0
    x"00",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D8
    x"00",x"00",x"00",x"04",x"0A",x"04",x"00",x"00", -- 0x01E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
    x"00",x"00",x"00",x"04",x"0A",x"08",x"1C",x"08", -- 0x01F0
    x"08",x"28",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0208
    x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"08", -- 0x0210
    x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0218
    x"00",x"00",x"00",x"14",x"14",x"14",x"00",x"00", -- 0x0220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0228
    x"00",x"00",x"00",x"14",x"14",x"3E",x"14",x"3E", -- 0x0230
    x"14",x"14",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0238
    x"00",x"00",x"00",x"08",x"1E",x"28",x"1C",x"0A", -- 0x0240
    x"3C",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0248
    x"00",x"00",x"00",x"32",x"32",x"04",x"08",x"10", -- 0x0250
    x"26",x"26",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0258
    x"00",x"00",x"00",x"10",x"28",x"28",x"10",x"2A", -- 0x0260
    x"24",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
    x"00",x"00",x"00",x"08",x"08",x"10",x"00",x"00", -- 0x0270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0278
    x"00",x"00",x"00",x"08",x"10",x"20",x"20",x"20", -- 0x0280
    x"10",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
    x"00",x"00",x"00",x"08",x"04",x"02",x"02",x"02", -- 0x0290
    x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0298
    x"00",x"00",x"00",x"00",x"08",x"2A",x"1C",x"1C", -- 0x02A0
    x"2A",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
    x"00",x"00",x"00",x"00",x"08",x"08",x"3E",x"08", -- 0x02B0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C0
    x"08",x"08",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x02C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"00", -- 0x02D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E0
    x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E8
    x"00",x"00",x"00",x"00",x"02",x"04",x"08",x"10", -- 0x02F0
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"00",x"00",x"00",x"1C",x"22",x"26",x"2A",x"32", -- 0x0300
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0308
    x"00",x"00",x"00",x"08",x"18",x"08",x"08",x"08", -- 0x0310
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0318
    x"00",x"00",x"00",x"1C",x"22",x"02",x"1C",x"20", -- 0x0320
    x"20",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0328
    x"00",x"00",x"00",x"1C",x"22",x"02",x"04",x"02", -- 0x0330
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0338
    x"00",x"00",x"00",x"04",x"0C",x"14",x"24",x"3E", -- 0x0340
    x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0348
    x"00",x"00",x"00",x"3E",x"20",x"3C",x"02",x"02", -- 0x0350
    x"02",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0358
    x"00",x"00",x"00",x"1C",x"20",x"20",x"3C",x"22", -- 0x0360
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0368
    x"00",x"00",x"00",x"3E",x"02",x"04",x"08",x"10", -- 0x0370
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0378
    x"00",x"00",x"00",x"1C",x"22",x"22",x"1C",x"22", -- 0x0380
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0388
    x"00",x"00",x"00",x"1C",x"22",x"22",x"1E",x"02", -- 0x0390
    x"02",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00", -- 0x03A0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
    x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00", -- 0x03B0
    x"08",x"08",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"04",x"08",x"10",x"20",x"10", -- 0x03C0
    x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"00",x"00",x"00",x"3E",x"00",x"3E", -- 0x03D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"00",x"00",x"00",x"10",x"08",x"04",x"02",x"04", -- 0x03E0
    x"08",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
    x"00",x"00",x"00",x"1C",x"22",x"02",x"04",x"08", -- 0x03F0
    x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
    x"00",x"00",x"00",x"1C",x"22",x"02",x"1A",x"2A", -- 0x0400
    x"2A",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0408
    x"00",x"00",x"00",x"08",x"14",x"22",x"22",x"3E", -- 0x0410
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0418
    x"00",x"00",x"00",x"3C",x"12",x"12",x"1C",x"12", -- 0x0420
    x"12",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0428
    x"00",x"00",x"00",x"1C",x"22",x"20",x"20",x"20", -- 0x0430
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
    x"00",x"00",x"00",x"3C",x"12",x"12",x"12",x"12", -- 0x0440
    x"12",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0448
    x"00",x"00",x"00",x"3E",x"20",x"20",x"3C",x"20", -- 0x0450
    x"20",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0458
    x"00",x"00",x"00",x"3E",x"20",x"20",x"3C",x"20", -- 0x0460
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0468
    x"00",x"00",x"00",x"1E",x"20",x"20",x"26",x"22", -- 0x0470
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0478
    x"00",x"00",x"00",x"22",x"22",x"22",x"3E",x"22", -- 0x0480
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0488
    x"00",x"00",x"00",x"1C",x"08",x"08",x"08",x"08", -- 0x0490
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0498
    x"00",x"00",x"00",x"02",x"02",x"02",x"02",x"22", -- 0x04A0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04A8
    x"00",x"00",x"00",x"22",x"24",x"28",x"30",x"28", -- 0x04B0
    x"24",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B8
    x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20", -- 0x04C0
    x"20",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04C8
    x"00",x"00",x"00",x"22",x"36",x"2A",x"2A",x"22", -- 0x04D0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04D8
    x"00",x"00",x"00",x"22",x"32",x"2A",x"26",x"22", -- 0x04E0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E8
    x"00",x"00",x"00",x"1C",x"22",x"22",x"22",x"22", -- 0x04F0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F8
    x"00",x"00",x"00",x"3C",x"22",x"22",x"3C",x"20", -- 0x0500
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0508
    x"00",x"00",x"00",x"1C",x"22",x"22",x"22",x"2A", -- 0x0510
    x"24",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0518
    x"00",x"00",x"00",x"3C",x"22",x"22",x"3C",x"28", -- 0x0520
    x"24",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0528
    x"00",x"00",x"00",x"1C",x"22",x"10",x"08",x"04", -- 0x0530
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0538
    x"00",x"00",x"00",x"3E",x"08",x"08",x"08",x"08", -- 0x0540
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0548
    x"00",x"00",x"00",x"22",x"22",x"22",x"22",x"22", -- 0x0550
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0558
    x"00",x"00",x"00",x"22",x"22",x"22",x"14",x"14", -- 0x0560
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0568
    x"00",x"00",x"00",x"22",x"22",x"22",x"2A",x"2A", -- 0x0570
    x"36",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0578
    x"00",x"00",x"00",x"22",x"22",x"14",x"08",x"14", -- 0x0580
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0588
    x"00",x"00",x"00",x"22",x"22",x"14",x"08",x"08", -- 0x0590
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0598
    x"00",x"00",x"00",x"3E",x"02",x"04",x"08",x"10", -- 0x05A0
    x"20",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A8
    x"00",x"00",x"00",x"38",x"20",x"20",x"20",x"20", -- 0x05B0
    x"20",x"38",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B8
    x"00",x"00",x"00",x"20",x"20",x"10",x"08",x"04", -- 0x05C0
    x"02",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C8
    x"00",x"00",x"00",x"0E",x"02",x"02",x"02",x"02", -- 0x05D0
    x"02",x"0E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D8
    x"00",x"00",x"00",x"08",x"1C",x"2A",x"08",x"08", -- 0x05E0
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E8
    x"00",x"00",x"00",x"00",x"08",x"10",x"3E",x"10", -- 0x05F0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F8
    x"00",x"00",x"00",x"08",x"14",x"22",x"00",x"00", -- 0x0600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0608
    x"00",x"00",x"00",x"00",x"00",x"1C",x"02",x"1E", -- 0x0610
    x"22",x"1E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0618
    x"00",x"00",x"00",x"20",x"20",x"2C",x"32",x"22", -- 0x0620
    x"32",x"2C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0628
    x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"20", -- 0x0630
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0638
    x"00",x"00",x"00",x"02",x"02",x"1A",x"26",x"22", -- 0x0640
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0648
    x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"3E", -- 0x0650
    x"20",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0658
    x"00",x"00",x"00",x"04",x"0A",x"08",x"1C",x"08", -- 0x0660
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0668
    x"00",x"00",x"00",x"00",x"00",x"1A",x"26",x"26", -- 0x0670
    x"1A",x"02",x"1C",x"00",x"00",x"00",x"00",x"00", -- 0x0678
    x"00",x"00",x"00",x"20",x"20",x"2C",x"32",x"22", -- 0x0680
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0688
    x"00",x"00",x"00",x"00",x"08",x"00",x"18",x"08", -- 0x0690
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0698
    x"00",x"00",x"00",x"00",x"02",x"00",x"02",x"02", -- 0x06A0
    x"02",x"22",x"1C",x"00",x"00",x"00",x"00",x"00", -- 0x06A8
    x"00",x"00",x"00",x"20",x"20",x"24",x"28",x"30", -- 0x06B0
    x"28",x"24",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06B8
    x"00",x"00",x"00",x"18",x"08",x"08",x"08",x"08", -- 0x06C0
    x"08",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C8
    x"00",x"00",x"00",x"00",x"00",x"14",x"2A",x"2A", -- 0x06D0
    x"2A",x"2A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D8
    x"00",x"00",x"00",x"00",x"00",x"2C",x"32",x"22", -- 0x06E0
    x"22",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06E8
    x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"22", -- 0x06F0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06F8
    x"00",x"00",x"00",x"00",x"00",x"2C",x"32",x"32", -- 0x0700
    x"2C",x"20",x"20",x"00",x"00",x"00",x"00",x"00", -- 0x0708
    x"00",x"00",x"00",x"00",x"00",x"1A",x"26",x"26", -- 0x0710
    x"1A",x"02",x"02",x"00",x"00",x"00",x"00",x"00", -- 0x0718
    x"00",x"00",x"00",x"00",x"00",x"2C",x"32",x"20", -- 0x0720
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0728
    x"00",x"00",x"00",x"00",x"00",x"1E",x"20",x"1C", -- 0x0730
    x"02",x"3C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0738
    x"00",x"00",x"00",x"10",x"10",x"38",x"10",x"10", -- 0x0740
    x"12",x"0C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0748
    x"00",x"00",x"00",x"00",x"00",x"22",x"22",x"22", -- 0x0750
    x"26",x"1A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0758
    x"00",x"00",x"00",x"00",x"00",x"22",x"22",x"22", -- 0x0760
    x"14",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0768
    x"00",x"00",x"00",x"00",x"00",x"22",x"2A",x"2A", -- 0x0770
    x"14",x"14",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
    x"00",x"00",x"00",x"00",x"00",x"22",x"14",x"08", -- 0x0780
    x"14",x"22",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0788
    x"00",x"00",x"00",x"00",x"00",x"22",x"22",x"22", -- 0x0790
    x"1E",x"02",x"1C",x"00",x"00",x"00",x"00",x"00", -- 0x0798
    x"00",x"00",x"00",x"00",x"00",x"3E",x"04",x"08", -- 0x07A0
    x"10",x"3E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A8
    x"00",x"00",x"00",x"08",x"10",x"10",x"20",x"10", -- 0x07B0
    x"10",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B8
    x"00",x"00",x"00",x"08",x"08",x"08",x"00",x"08", -- 0x07C0
    x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
    x"00",x"00",x"00",x"08",x"04",x"04",x"02",x"04", -- 0x07D0
    x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D8
    x"00",x"00",x"00",x"10",x"2A",x"04",x"00",x"00", -- 0x07E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F0
    x"00",x"3E",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x07F8
	
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
	    DATA_R <= RAM(to_integer(unsigned(ADDR_R)));
		if WE = '1' then
			RAM(to_integer(unsigned(ADDR_W))) <= DATA_W;
		end if;
  end process;
end RTL;
